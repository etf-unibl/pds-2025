-----------------------------------------------------------------------------
-- Faculty of Electrical Engineering
-- PDS 2025
-- https://github.com/etf-unibl/pds-2025/
-----------------------------------------------------------------------------
--
-- unit name:     single_digit_bcd_adder
--
-- description:
--
--   This file implements single digit BCD adder
--
-----------------------------------------------------------------------------
-- Copyright (c) 2025 Faculty of Electrical Engineering
-----------------------------------------------------------------------------
-- The MIT License
-----------------------------------------------------------------------------
-- Copyright 2025 Faculty of Electrical Engineering
--
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the "Software"),
-- to deal in the Software without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Software, and to permit persons to whom
-- the Software is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
-- THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity single_digit_bcd_adder is
	port (
	A_i   : in std_logic_vector(3 downto 0);
	B_i   : in std_logic_vector(3 downto 0);
	CARRY_i : in std_logic;
	SUM_o : out std_logic_vector(3 downto 0);
	CARRY_o : out std_logic
);
end single_digit_bcd_adder;

architecture single_digit_bcd_adder_arch of single_digit_bcd_adder is
begin
process(A_i, B_i, CARRY_i)
	variable temp : unsigned(4 downto 0);
begin
	temp := unsigned('0'&A_i) + unsigned('0'&B_i) + ("0000"&CARRY_i);
	if(temp > 9) then
		CARRY_o <= '1';
		SUM_o <= std_logic_vector(resize((temp + "00110"),4));
	else
		CARRY_o <= '0';
		SUM_o <= std_logic_vector(resize(temp, 4));
	end if;
end process;
end architecture;
