library ieee;
use ieee.std_logic_1164.all;

entity test is
end entity test;

architecture rtl of test is
begin
	--Prazna arhitektura
end architecture rtl;