-- File: test.vhd
-- Minimalni VHDL dizajn: entitet sa praznom arhitekturom

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity test is
end entity test;

architecture empty of test is
begin
    -- Prazna arhitektura
end architecture empty;