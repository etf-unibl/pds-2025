library ieee;

use ieee.std_logic_1164.all;

entity test is


	
end test;

architecture test_arch of test is
	

end test_arch;