library ieee;

use ieee.std_logic_1164.all;

entity test is	

end entity test;

architecture test_arch of test is
begin	
end architecture test_arch;