library IEEE;
use IEE.STD_LOGIC_1164.ALL;

entity test is 
end entity test;

architecture arch of test is
begin
	--empty 
end architecture arch;