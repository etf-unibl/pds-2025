library ieee;
use ieee.std_logic_1164.all;

entity d_ff_tb is 
end entity d_ff_tb;

architecture rtl of d_ff_tb is 
begin
    -- empty
end architecture rtl;
